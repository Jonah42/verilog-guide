`timescale 1ns / 1ps

// Jonah Meggs 2022
// Jonah's Guide to Verilog Chapter 1 - minimal.v
// The simplest example of Verilog I can think of

module minimal(
	output o
    );

assign o = 1;

endmodule
