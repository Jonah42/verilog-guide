`timescale 1ns / 1ps

// Jonah Meggs 2022
// Jonah's Guide to Verilog Chapter 1 - minimal2.v
// Adding input to minimal.v

module minimal2(
	input i,
	output o
    );

assign o = i;

endmodule
